class c_184_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_184_4;
    c_184_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01zz11x10x01xz1x101xz100z0x0000xzzzzxxzxzxxzxzxzxxzxxxzxxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
