class c_182_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_182_1;
    c_182_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xzx0xx011xxx10x10x00xx11x1zzz0zzxxxxzzxxxxzxzzzzzxzxzxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
