class c_49_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_49_4;
    c_49_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz0xxz11z1111x0xzx0011zx0xx0xx0zzzzxxzzxzzxzzzxxzxzzzxzzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
