`define SMC_MCPER_ADDR       7'h00
`define SMC_MCCTL1_ADDR       7'h02
`define SMC_MCCTL0_ADDR       7'h03
`define SMC_MCCC3_ADDR       7'h10
`define SMC_MCCC2_ADDR       7'h11
`define SMC_MCCC1_ADDR       7'h12
`define SMC_MCCC0_ADDR       7'h13
`define SMC_MCCC7_ADDR       7'h14
`define SMC_MCCC6_ADDR       7'h15
`define SMC_MCCC5_ADDR       7'h16
`define SMC_MCCC4_ADDR       7'h17
`define SMC_MCCC11_ADDR       7'h18
`define SMC_MCCC10_ADDR       7'h19
`define SMC_MCCC9_ADDR       7'h1A
`define SMC_MCCC8_ADDR       7'h1B
`define SMC_MCDC1_ADDR       7'h20
`define SMC_MCDC0_ADDR       7'h22
`define SMC_MCDC3_ADDR       7'h24
`define SMC_MCDC2_ADDR       7'h26
`define SMC_MCDC5_ADDR       7'h28
`define SMC_MCDC4_ADDR       7'h2A
`define SMC_MCDC7_ADDR       7'h2C
`define SMC_MCDC6_ADDR       7'h2E
`define SMC_MCDC9_ADDR       7'h30
`define SMC_MCDC8_ADDR       7'h32
`define SMC_MCDC11_ADDR       7'h34
`define SMC_MCDC10_ADDR       7'h36
