class c_192_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_192_1;
    c_192_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zzzzz1z0zzzxxx00zxx1zx01100z00xzxzzxzzxzzzzzzzxzzxxxxxzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
