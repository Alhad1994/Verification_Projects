class c_137_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_137_1;
    c_137_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z10xx010x0100z0x110x1z0xzx111zxxxxzzzxzzxxxxzzxxzxxxzzxxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
