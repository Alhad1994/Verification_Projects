`include "./../seq/base_seq.sv"
`include "./../seq/reg_seq.sv"
`include "./../seq/per_seq.sv"
`include "./../seq/smc_seq.sv"
`include "./../uvc/smc_sequencer.sv"
`include "./../uvc/smc_driver.sv"
`include "./../uvc/smc_monitor.sv"
`include "./../uvc/smc_scoreboard.sv"
`include "./../uvc/smc_agent.sv"
`include "./../uvc/smc_env.sv"
`include "./../test/reg_test.sv"
`include "./../test/per_test.sv"
`include "./../test/smc_test.sv"
