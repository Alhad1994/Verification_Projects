class c_54_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_54_4;
    c_54_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xzzz1xz000z0xzxxx00z00xz1zzzx0xzxxzxxzzxxzxxzzzxxxzxzzzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
