class c_197_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_197_4;
    c_197_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzzx1xxzz0z1011100xz01011xzx00xzzzxzzxzxzzxzxzxzzzxxxzzxzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
