class c_178_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_178_4;
    c_178_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx0x000zx0xz111xxzxx00xz0x0xz11xxxzxxzzzzxxzxzzzzxzxxzzzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
