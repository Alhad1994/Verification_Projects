class c_142_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_142_4;
    c_142_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001zz0x000x01xz000zz10x101x01111zxzzzzzzzzzzzxzxxxzxzxzxxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
