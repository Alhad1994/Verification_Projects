class c_156_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_156_4;
    c_156_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx1z1xx01101x0x0z10x11xzzzz0zx1zxzxzxzzxxxxxxxxzzxzzzzzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
