class c_49_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_49_1;
    c_49_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zx0xx1zz1010x0z0zxx10x0z0zx0zzxzzzzxxxxzxzxxzxzzzxzzzxzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
