class c_128_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_128_1;
    c_128_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x100101xx1z010xx01x0xzz1011z0zxxxxzxzxzzxxzzzzxxxxzzxxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
