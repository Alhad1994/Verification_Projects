class c_181_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_181_4;
    c_181_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zz1z1xxzzzxx0001xz1zx0z0x0z1zzzxzxzxxxxzxzxzzzxzzxxzxzzxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
