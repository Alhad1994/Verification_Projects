class c_97_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_97_4;
    c_97_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz1xzzx10x11zx1xx0x1xxzzx11x01zxxxxzzxxxxxxxzxxzxxxzxxzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
