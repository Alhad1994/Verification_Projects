class c_24_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_24_1;
    c_24_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z101z0zzx01xxx1z1z000z0xz1zzx1zzxzzxzxxxxxxxxxxzxzzxxxzxxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
