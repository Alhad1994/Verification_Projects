class c_138_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_138_4;
    c_138_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz101zz0zx01zx11z1011110zzx0xxxzzxzxxxzzzxxxzxxxxxzzxxxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
