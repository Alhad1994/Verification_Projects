class c_102_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_102_1;
    c_102_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z011xz1zx11111zx01z00x0x0zzzz0zzxxxxxzzzzxzxzzxzxzxzzxxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
