class c_60_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_60_1;
    c_60_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0110zz01xz0xzx1xzxxx1z10zx0xxxzxzxzzzxxzxzxzxzxxxzzzxzzxxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
