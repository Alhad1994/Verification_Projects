class c_20_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_20_1;
    c_20_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01zzzz1zxzx1z110xzxz1x10xz1xzzxxzxxzzxxzxzxzxxxzzxxzxzxzxxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
