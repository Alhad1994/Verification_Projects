class c_97_1;
    rand bit[25:0] clk_freq; // rand_mode = ON 

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_97_1;
    c_97_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz01x00x11xx1x1111xxz001z00zx00zxxxxzxxxxzxzzxzzzxzzzzxzxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
