class c_98_4;
    bit[25:0] clk_freq = 26'hf4240;

    constraint freq_this    // (constraint_mode = ON) (./../seq/uart_tr.sv:27)
    {
       ((clk_freq[25]) == ((clk_freq[25]) + 5));
    }
endclass

program p_98_4;
    c_98_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100z001zx1zzxxz0xx0011xx0x1zzxzzzxzxzxzzxzxzzzzzxxxzzxxzxxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
